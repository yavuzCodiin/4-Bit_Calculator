library IEEE; 
use IEEE.STD_LOGIC_1164.ALL; 
use IEEE.STD_LOGIC_ARITH.ALL; 
use IEEE.STD_LOGIC_UNSIGNED.ALL; 

ENTITY MUXTWOTONE IS
PORT (
		 A0 : IN STD_LOGIC_VECTOR (3 DOWNTO 0); 
		 A1  : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		 S  : IN STD_LOGIC;
		 OUTPUT : OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
END MUXTWOTONE;
ARCHITECTURE Behavior OF MUXTWOTONE IS	
BEGIN
	WITH S SELECT
		    OUTPUT <= 	A0 WHEN '0',
						A1 WHEN  OTHERS;
END Behavior;
