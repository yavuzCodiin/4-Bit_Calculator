library IEEE; 
use IEEE.STD_LOGIC_1164.ALL; 
use IEEE.STD_LOGIC_ARITH.ALL; 
use IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY EIGHTTOONEMUX IS
	PORT (
		 RA : IN STD_LOGIC_VECTOR (3 DOWNTO 0); 
		 LLS  : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		 LRS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		 ARS  : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		 RB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		 RBINV  : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		 DIN  : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		 DIINV : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		 IN_SELECT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		 OUTPUT : OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
END EIGHTTOONEMUX;
ARCHITECTURE Behavior OF EIGHTTOONEMUX IS	
BEGIN
	WITH IN_SELECT SELECT
		    OUTPUT <= 	
					RA WHEN "000", 
					LLS WHEN "001", 
					LRS WHEN "010", 
					ARS WHEN "011", 
            		RB WHEN "100", 
             		RBINV WHEN "101", 
            		DIN WHEN "110",
             		DIINV WHEN OTHERS;
END Behavior;
